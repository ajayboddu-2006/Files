magic
tech min2
timestamp 1712917271
<< nwell >>
rect -7 -4 11 11
<< nsubstratencontact >>
rect -9 -14 -6 -11
<< polysilicon >>
rect -13 -14 -10 -11
<< end >>
