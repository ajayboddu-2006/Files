\m5_TLV_version 1d: tl-x.org
\m5
\SV
   m5_makerchip_module   
\TLV
  //Logic Gates
  $out1 = $in1 & $in2;
  $out2 = $in1 | $in2;
  $out3 = ~$in1;
  $out4 = !($in1 & $in2);
  $out5 = !($in1 | $in2);
  $out6 = !($in1 ^ $in2);
  $out7 = $in1 ^ $in2;
  
\SV
   endmodule
